module TestBenchQ2_1;
	reg [31:0] Num_1;
	reg [31:0] Num_2;
	reg [31:0] Num_3;
	reg [31:0] Num_4;
	reg [31:0] Num_5;
	reg [31:0] Num_6;
	reg [31:0] Num_7;
	reg [31:0] Num_8;
	reg [31:0] Num_9;
	reg [31:0] Num_10;
	reg [31:0] Num_11;
	reg [31:0] Num_12;
	reg [31:0] Num_13;
	reg [31:0] Num_14;
	reg [31:0] Num_15;
	reg [31:0] Num_16;
	reg [31:0] Target_Num;
	reg Clock = 0;
	reg Reset;
	wire [3:0] Out_4;
	
	Correlation_32 module_test_Q2_1(Num_1, Num_2, Num_3, Num_4, Num_5, Num_6, Num_7, Num_8, Num_9, Num_10, Num_11, Num_12, Num_13, Num_14, Num_15, Num_16, Target_Num, Clock, Reset, Out_4);
	always forever begin #10 Clock = ~Clock;
	end	
	initial
	begin
		Reset = 0;
		#5;
		Reset = 1;
		#5;
		Reset = 0;
		Target_Num = 60;
		$display("Target_Num = %b",Target_Num);
		Num_1 = $dist_normal($time, 100, 20);
		Num_2 = $dist_normal($time, 200, 20);
		Num_3 = $dist_normal($time, 300, 20);
		Num_4 = $dist_normal($time, 400, 20);
		Num_5 = $dist_normal($time, 50, 20);
		Num_6 = $dist_normal($time, 60, 20);
		Num_7 = $dist_normal($time, 70, 20);
		Num_8 = $dist_normal($time, 80, 20);
		Num_9 = $random();
		Num_10 = $random();
		Num_11 = $random();
		Num_12 = $random();
		Num_13 = $random();
		Num_14 = $random();
		Num_15 = $random();
		Num_16 = $random();
		#20;
		$display("RESET IS %s" ,Reset ? "ON" : "OFF");
		$display("Num_1 = %b",Num_1);
		$display("Num_2 = %b",Num_2);
		$display("Num_3 = %b",Num_3);
		$display("Num_4 = %b",Num_4);
		$display("Num_5 = %b",Num_5);
		$display("Num_6 = %b",Num_6);
		$display("Num_7 = %b",Num_7);
		$display("Num_8 = %b",Num_8);
		$display("Num_9 = %b",Num_9);
		$display("Num_10 = %b",Num_10);
		$display("Num_11 = %b",Num_11);
		$display("Num_12 = %b",Num_12);
		$display("Num_13 = %b",Num_13);
		$display("Num_14 = %b",Num_14);
		$display("Num_15 = %b",Num_15);
		$display("Num_16 = %b",Num_16);
		$display("Congratulation Player %d! You are the winner!", Out_4);
		Target_Num = 30;
		$display("Target_Num = %b",Target_Num);
		Num_1 = $random();
		Num_2 = $random();
		Num_3 = $random();
		Num_4 = $random();
		Num_5 = $random();
		Num_6 = $random();
		Num_7 = $random();
		Num_8 = $random();
		Num_9 = $dist_normal($time, 80, 20);
		Num_10 = $dist_normal($time, 70, 20);
		Num_11 = $dist_normal($time, 60, 20);
		Num_12 = $dist_normal($time, 50, 20);
		Num_13 = $dist_normal($time, 400, 20);
		Num_14 = $dist_normal($time, 300, 20);
		Num_15 = $dist_normal($time, 200, 20);
		Num_16 = $dist_normal($time, 100, 20);
		#20;
		$display("RESET IS %s" ,Reset? "ON" : "OFF");
		$display("Num_1 = %b",Num_1);
		$display("Num_2 = %b",Num_2);
		$display("Num_3 = %b",Num_3);
		$display("Num_4 = %b",Num_4);
		$display("Num_5 = %b",Num_5);
		$display("Num_6 = %b",Num_6);
		$display("Num_7 = %b",Num_7);
		$display("Num_8 = %b",Num_8);
		$display("Num_9 = %b",Num_9);
		$display("Num_10 = %b",Num_10);
		$display("Num_11 = %b",Num_11);
		$display("Num_12 = %b",Num_12);
		$display("Num_13 = %b",Num_13);
		$display("Num_14 = %b",Num_14);
		$display("Num_15 = %b",Num_15);
		$display("Num_16 = %b",Num_16);
		$display("Congratulation Player %d! You are the winner!", Out_4);
		#100;
		Reset = 1;
	end     
endmodule