module SixteenToOneMultiplexerWithThirtyTwoBitLength
(
input_1,
input_2,
input_3,
input_4,
input_5,
input_6,
input_7,
input_8,
input_9,
input_10,
input_11,
input_12,
input_13,
input_14,
input_15,
input_16,
select,
output_1
);
input [31:0] input_1;
input [31:0] input_2;
input [31:0] input_3;
input [31:0] input_4;
input [31:0] input_5;
input [31:0] input_6;
input [31:0] input_7;
input [31:0] input_8;
input [31:0] input_9;
input [31:0] input_10;
input [31:0] input_11;
input [31:0] input_12;
input [31:0] input_13;
input [31:0] input_14;
input [31:0] input_15;
input [31:0] input_16;
input [4:0] select;
output [31:0] output_1;
wire [31:0] WIRE_1[3:0];
wire [31:0] WIRE_2[3:0];
wire [1:0] WIRE_select;
assign WIRE_select[0] = select[4];
assign WIRE_select[1] = 1'b0;
assign WIRE_2[2] = 0;
assign WIRE_2[1] = 0;
assign WIRE_2[0] = 0;
FourToOneMultiplexerWithThirtyTwoBitLength Test_0(input_1, input_2, input_3, input_4, select[1:0], WIRE_1[3]);
FourToOneMultiplexerWithThirtyTwoBitLength Test_1(input_5, input_6, input_7, input_8, select[1:0], WIRE_1[2]);
FourToOneMultiplexerWithThirtyTwoBitLength Test_2(input_9, input_10, input_11, input_12, select[1:0], WIRE_1[1]);
FourToOneMultiplexerWithThirtyTwoBitLength Test_3(input_13, input_14, input_15, input_16, select[1:0], WIRE_1[0]);
FourToOneMultiplexerWithThirtyTwoBitLength Test_4(WIRE_1[3], WIRE_1[2], WIRE_1[1], WIRE_1[0], select[3:2], WIRE_2[3]);
FourToOneMultiplexerWithThirtyTwoBitLength Test_5(WIRE_2[3], WIRE_2[2], WIRE_2[1], WIRE_2[0], WIRE_select, output_1);
endmodule